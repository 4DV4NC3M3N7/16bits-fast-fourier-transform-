
module FFT (
	clk_clk);	

	input		clk_clk;
endmodule
